//-------------------------------------------------------------------------
//    Color_Mapper.sv                                                    --
//    Stephen Kempf                                                      --
//    3-1-06                                                             --
//                                                                       --
//    Modified by David Kesler  07-16-2008                               --
//    Translated by Joe Meng    07-07-2013                               --
//                                                                       --
//    Fall 2014 Distribution                                             --
//                                                                       --
//    For use with ECE 385 Lab 7                                         --
//    University of Illinois ECE Department                              --
//-------------------------------------------------------------------------

module  color_mapper ( input        [9:0] user1X, user1Y, bomb1X, bomb1Y, bomb1S, user1S,
							  input 			[9:0] user2X, user2Y, bomb2X, bomb2Y, bomb2S, user2S,
							  input        [9:0] wall1X, wall1Y, wall1S,
							  input		   [9:0] DrawX, DrawY,
							  input			Clk, blank,
							  
                       output logic [7:0]  Red, Green, Blue);
							  
  logic user1_on, bomb1_on, user2_on, bomb2_on;
  logic wall1_on;

	 logic [7:0] TR, TG, TB;
   logic [23:0] temp_data;
/* 
     New Ball: Generates (pixelated) circle by using the standard circle formula.  Note that while 
     this single line is quite powerful descriptively, it causes the synthesis tool to use up three
     of the 12 available multipliers on the chip!  Since the multiplicants are required to be signed,
	  we have to first cast them from logic to int (signed by default) before they are multiplied). 
*/
	  
    logic [9:0] user1DistX, user1DistY;
	 
	 int user1Size, bomb1DistX, bomb1DistY, bomb1Size;
	 int user2DistX, user2DistY, user2Size, bomb2DistX, bomb2DistY, bomb2Size;
	 int wall1DistX, wall1DistY, wall1Size;
	 
	 assign wall1Size = wall1S;
	 assign wall1DistX = DrawX - wall1X;
    assign wall1DistY = DrawY - wall1Y;
	 
    assign user1Size = user1S;	 
  	 assign user1DistX = DrawX - user1X; //(x-h) 
    assign user1DistY = DrawY - user1Y;
	 
	 assign bomb1DistX = DrawX - bomb1X;
    assign bomb1DistY = DrawY - bomb1Y;
    assign bomb1Size = bomb1S;
	 
	 assign user2DistX = DrawX - user2X;
    assign user2DistY = DrawY - user2Y;
    assign user2Size = user2S;
	 

	 assign bomb2DistX = DrawX - bomb2X;
    assign bomb2DistY = DrawY - bomb2Y;
    assign bomb2Size = bomb2S;
 
	 
logic [18:0] addr;
logic [3:0] rom_addr;
	 
assign addr = user1DistX + (16 * user1DistY);

background_ram sprite1(  .read_address(addr),
									.Clk(Clk),
									.data_Out(temp_data));	
//map ram
//bomb ram
					

always_ff @(posedge Clk) 
	begin
		TR [7:0]	<= temp_data[23:16];
		TG [7:0] <= temp_data[15:8];
		TB [7:0] <= temp_data[7:0];
		
	end

    always_comb
    begin
			//User 1 display
        if ((user1DistX <= 10'd16 && user1DistY <= 10'd23) && ((user1DistX >= 10'd0 && user1DistY >= 10'd0))) 
				begin
					user1_on = 1'b1;
				end
				
			else 
			 begin
					user1_on = 1'b0;
			 end

			
				//Bomb 1 Display
		  if ( ( bomb1DistX*bomb1DistX + bomb1DistY*bomb1DistY) <= (bomb1Size * bomb1Size) ) 
			begin
            bomb1_on = 1'b1;
			end
			
		  else 
			begin
				bomb1_on = 1'b0;
			end
			
			// User 2 Display
			if ( ( user2DistX*user2DistX + user2DistY*user2DistY) <= (user2Size * user2Size) ) 
			begin
            user2_on = 1'b1;
			end
			
		  else 
			begin
				user2_on = 1'b0;
			end
		
			//Bomb 2 Display
		  if ( ( bomb2DistX*bomb2DistX + bomb2DistY*bomb2DistY) <= (bomb2Size * bomb2Size) ) 
			begin
            bomb2_on = 1'b1;
			end
			
		  else 
			begin
				bomb2_on = 1'b0;
			end
			
        //  Wall Display
		  
        if ((wall1DistX < wall1S && wall1DistY < wall1S) && ((wall1DistX >= 10'd0 && wall1DistY >= 10'd0)))
			begin
            wall1_on = 1'b1;
			end
			
		  else 
			begin
				wall1_on = 1'b0;
			end
		 
		  
end


 always_ff @ (posedge Clk)
    begin:RGB_Display
       
	  if(blank)
		begin

		 if ((user1_on == 1'b1)) 
		  begin
			
				
				Red <= TR;
				Green <= TG;
				Blue <= TB;
				
			end 
		  
		  else if ((bomb1_on == 1'b1))
		  begin
				Red = 8'h00;
				Green = 8'hff;
				Blue = 8'h00;

			end
			
		  else if ((bomb2_on == 1'b1))
		  begin
				Red = 8'h00;
				Green = 8'hff;
				Blue = 8'h00;
		  
		  end
		  
		  else if ((user2_on == 1'b1)) 
        begin 
            Red = 8'h00;
            Green = 8'h00;
            Blue = 8'hFF;

        end 
		  
		  else if ((wall1_on == 1'b1)) 
        begin 
            Red = 8'hFF;
            Green = 8'hFF;
            Blue = 8'hFF;

        end 
		  
		  else
        begin 
            Red = 8'h00; 
            Green = 8'h00;
            Blue = 8'h7f - DrawX[9:3];
        end 
		  
		 end
		  
        else
        begin 
            Red = 8'h00; 
            Green = 8'h00;
            Blue = 8'h00;

        end 
		
    end 
    
endmodule 